LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY delta_example_tb IS
END delta_example_tb;

ARCHITECTURE tb OF delta_example_tb IS
    SIGNAL S : INTEGER := 0;
BEGIN

    stim_pro : PROCESS
        VARIABLE V : INTEGER := 0;

    BEGIN
        REPORT "=== Inicio del proceso ===";

        -- Primera asignaci�n
        V := 1;
        S <= 1;
        REPORT "Delta 1: V=" & INTEGER'IMAGE(V) & ", S=" & INTEGER'IMAGE(S);

        -- Segunda asignaci�n
        V := 2;
        S <= 2;
        REPORT "Delta 2: V=" & INTEGER'IMAGE(V) & ", S=" & INTEGER'IMAGE(S);

        -- Tercera asignaci�n
        V := 3;
        S <= 3;
        REPORT "Delta 3: V=" & INTEGER'IMAGE(V) & ", S=" & INTEGER'IMAGE(S);

        -- Ahora esperamos una actualizaci�n de se�ales
        WAIT FOR 0 ns;

        REPORT "Despu�s de WAIT FOR de 0 ns: V=" & INTEGER'IMAGE(V) & ", S=" & INTEGER'IMAGE(S);

        WAIT; -- Detener la simulaci�n

    END PROCESS;
END tb;